module test_inputs(
);